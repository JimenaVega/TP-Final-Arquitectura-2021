`timescale 1ns / 1ps

module TOP#(

    )
    (
        input                       i_clock,
        input                       i_reset
    );
    
    IF_stage IF_stage_1(.i_clock(),
                        .i_IF_branch(),
                        .i_IF_jump(),
                        .i_IF_pc_enable(),
                        .i_IF_pc_reset(),
                        .i_IF_read_enable(),
                        .i_IF_branch_address(),
                        .i_IF_jump_address(),
                        .o_IF_adder_result(),
                        .o_IF_new_instruction());
                        
    IF_ID_reg IF_ID_reg_1(.i_clock(),
                          .IF_adder_result(),
                          .IF_new_instruction(),
                          .ID_adder_result(),
                          .ID_new_instruction());
    
    ID_stage ID_stage_1(.i_ID_clock(),
                        .i_ID_reset(),
                        .i_ID_enable(),
                        .i_ID_inst(),
                        .i_ID_pc(),
                        .i_ID_write_data(),
                        .i_ID_write_reg(),
                        .i_ID_reg_write(),
                        .o_ID_reg_dest(),
                        .o_ID_alu_op(),
                        .o_ID_alu_src(),
                        .o_ID_mem_read(),
                        .o_ID_mem_write(),
                        .o_ID_branch(),
                        .o_ID_reg_write(),
                        .o_ID_mem_to_reg(),
                        .o_ID_jump(),
                        .o_ID_jump_address(),
                        .o_ID_data_a(),
                        .o_ID_data_b(),
                        .o_ID_immediate(),
                        .o_ID_rt(),
                        .o_ID_rd(),
                        .o_ID_pc());
                        
    ID_EX_reg ID_EX_reg_1(.i_clock(),
                          .ID_reg_write(),
                          .ID_mem_to_reg(),
                          .ID_mem_read(),
                          .ID_mem_write(),
                          .ID_branch(),
                          .ID_alu_src(),
                          .ID_reg_dst(),
                          .ID_alu_op(),
                          .ID_pc(),
                          .ID_data_a(),
                          .ID_data_b(),
                          .ID_immediate(),
                          .ID_rt(),
                          .ID_rd(),
                          .EX_reg_write(),
                          .EX_mem_to_reg(),
                          .EX_mem_read(),
                          .EX_mem_write(),
                          .EX_branch(),
                          .EX_alu_src(),
                          .EX_reg_dst(),
                          .EX_alu_op(),
                          .EX_pc(),
                          .EX_data_a(),
                          .EX_data_b(),
                          .EX_immediate(),
                          .EX_rt(),
                          .EX_rd());
    
    EX_stage EX_stage_1(.i_clock(),
                        .i_EX_reg_write(),
                        .i_EX_mem_to_reg(),
                        .i_EX_mem_read(),
                        .i_EX_mem_write(),
                        .i_EX_branch(),
                        .i_EX_alu_src(),
                        .i_EX_reg_dst(),
                        .i_EX_alu_op(),
                        .i_EX_pc(),
                        .i_EX_data_a(),
                        .i_EX_data_b(),
                        .i_EX_immediate(),
                        .i_EX_rt(),
                        .i_EX_rd(),
                        .o_EX_reg_write(),
                        .o_EX_mem_to_reg(),
                        .o_EX_mem_read(),
                        .o_EX_mem_write(),
                        .o_EX_branch(),
                        .o_EX_branch_address(),
                        .o_EX_zero(),
                        .o_EX_alu_result(),
                        .o_EX_data_a(),
                        .o_EX_selected_reg());
                        
    EX_MEM_reg EX_MEM_reg_1(.i_clock(),
                            .EX_reg_write(),
                            .EX_mem_to_reg(),
                            .EX_mem_read(),
                            .EX_mem_write(),
                            .EX_branch(),
                            .EX_branch_address(),
                            .EX_zero(),
                            .EX_alu_result(),
                            .EX_data_a(),
                            .EX_selected_reg(),
                            .MEM_reg_write(),
                            .MEM_mem_to_reg(),
                            .MEM_mem_read(),
                            .MEM_mem_write(),
                            .MEM_branch(),
                            .MEM_branch_address(),
                            .MEM_zero(),
                            .MEM_alu_result(),
                            .MEM_data_a(),
                            .MEM_selected_reg());
                
    MEM_stage MEM_stage_1(.i_clock(),
                          .i_reset(),
                          .i_MEM_reg_write(),
                          .i_MEM_mem_to_reg(),
                          .i_MEM_mem_read(),
                          .i_MEM_mem_write(),
                          .i_MEM_word_en(),
                          .i_MEM_halfword_en(),
                          .i_MEM_byte_en(),
                          .i_MEM_branch(),
                          .i_MEM_zero(),
                          .i_MEM_branch_addr(),
                          .i_MEM_alu_result(),
                          .i_MEM_write_data(),
                          .i_MEM_selected_reg(),
                          .o_MEM_mem_data(),
                          .o_MEM_selected_reg(),
                          .o_MEM_alu_result(),
                          .o_MEM_branch_address(),
                          .o_branch_zero(),
                          .o_MEM_reg_write(),
                          .o_MEM_mem_to_reg());
                         
    MEM_WB_reg MEM_WB_reg_1(.i_clock(),
                            .i_MEM_reg_write(),
                            .i_MEM_mem_to_reg(),
                            .i_MEM_mem_data(),
                            .i_MEM_alu_result(),
                            .i_MEM_selected_reg(),
                            .o_WB_reg_write(),
                            .o_WB_mem_to_reg(),
                            .o_WB_mem_data(),
                            .o_WB_alu_result(),
                            .o_WB_selected_reg());
                          
    WB_stage WB_stage_1(.i_WB_reg_write(),
                        .i_WB_mem_to_reg(),
                        .i_WB_mem_data(),
                        .i_WB_alu_result(),
                        .i_WB_selected_reg(),
                        .o_WB_reg_write(),
                        .o_WB_selected_data(),
                        .o_WB_selected_reg());

endmodule
